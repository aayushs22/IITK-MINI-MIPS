`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/09/2025 02:32:52 PM
// Design Name: 
// Module Name: inst_file
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instr_fetch(input [14:0] addr, output [31:0] instr);
    reg [31:0] instr_mem[31:0];

    initial begin
        //instr_mem[0] <= 32'b001111_00000_00001_0000000000000001;
        //instr_mem[1] <= 32'b100001_00010_00001_01000_00000000011;
	//instr_mem[2] <= 32'b011010_00010_00001_00000_00011000111;
        //instr_mem[0] <= 32'b010010_00000_00001_0000000000000011;
        //instr_mem[1] <= 32'h0bc12345;
        


instr_mem[0]  <= 32'b000001_00000_00001_0000000000000001;
instr_mem[1]  <= 32'b010000_00100_00001_0000000000010010;
instr_mem[2]  <= 32'b000010_00001_00010_00000_00000_000001;
instr_mem[3]  <= 32'b010100_00010_00000_0000000000010000;
instr_mem[4]  <= 32'b100001_00011_00010_01001_00000_000000;
instr_mem[5]  <= 32'b001110_01001_00101_0000000000000000;
instr_mem[6]  <= 32'b001110_01001_00110_0000000000000001;
instr_mem[7]  <= 32'b101100_00110_00101_00111_00000_000000;
instr_mem[8]  <= 32'b010000_00000_00111_0000000000001110;
instr_mem[9]  <= 32'b000001_00110_01000_0000000000000000;
instr_mem[10] <= 32'b000001_00101_00110_0000000000000000;
instr_mem[11] <= 32'b000001_01000_00101_0000000000000000;
instr_mem[12] <= 32'b001111_01001_00101_0000000000000000;
instr_mem[13] <= 32'b001111_01001_00110_0000000000000001;
instr_mem[14] <= 32'b000010_00010_00010_00000_00000_000001;
instr_mem[15] <= 32'b011000_00000000000_000000000000011;
instr_mem[16] <= 32'b000001_00001_00001_0000000000000001;
instr_mem[17] <= 32'b011000_00000000000_000000000000001;

    end

    assign instr = instr_mem[addr];
endmodule
